.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.064pF, R0=100ohm, Rn=16ohm, Icrit=0.1mA)
.model pjjmod jj(Rtype=1, Vg=2.8mV, Cap=0.064pF, R0=100ohm, Rn=16ohm, Icrit=0.1mA, PHI=PI)


** + -------------------- +
** |     HFQJTL           |
** + -------------------- +

.subckt jtl_squid   2       5 
L0 2 3 0.00001pH
L1 3 1 1.2pH
L2 3 4 1.2pH
B1 1 5 jjmod area=0.7440000000000001
R1 1 5 10.39ohm
B2 4 5 pjjmod area=0.7440000000000001
R2 4 5 10.39ohm
.ends

.subckt jtl_base        1       5       100
L1 1 2 0.684pH
L2 2 3 2.874pH
L3 3 4 5.748pH
L4 4 5 2.19pH
X1      jtl_squid       3       0
X2      jtl_squid       4       0
R1 2 100 25.01ohm
.ends


.subckt jtl_base8       1       9       100
X1      jtl_base        1       2       100
X2      jtl_base        2       3       100
X3      jtl_base        3       4       100
X4      jtl_base        4       5       100
X5      jtl_base        5       6       100
X6      jtl_base        6       7       100
X7      jtl_base        7       8       100
X8      jtl_base        8       9       100
.ends
** + -------------------- +



** + -------------------- +
** |     HFQJTL    test   |
** + -------------------- +
.subckt jtl_squid_test   2       5 
L0 2 3 0.00001pH
L1 3 1 1.2pH
L2 3 4 1.2pH
B1 1 5 jjmod area=0.7440000000000001
R1 1 5 10.39ohm
B2 4 5 pjjmod area=0.7440000000000001
R2 4 5 10.39ohm
.ends

.subckt jtl_base_test        1       5       100
L1 1 2 0.684pH
L2 2 3 2.874pH
L3 3 4 5.748pH
L4 4 5 2.19pH
X1      jtl_squid_test       3       0
X2      jtl_squid_test       4       0
R1 2 100 25.01ohm
.ends

.subckt jtl_base20       1       21       100
X1      jtl_base_test        1       2       100
X2      jtl_base_test        2       3       100
X3      jtl_base_test        3       4       100
X4      jtl_base_test        4       5       100
X5      jtl_base_test        5       6       100
X6      jtl_base_test        6       7       100
X7      jtl_base_test        7       8       100
X8      jtl_base_test        8       9       100
X9      jtl_base_test        9       10      100
X10     jtl_base_test       10       11      100
X11     jtl_base_test       11       12      100
X12     jtl_base_test       12       13      100
X13     jtl_base_test       13       14      100
X14     jtl_base_test       14       15      100
X15     jtl_base_test       15       16      100
X16     jtl_base_test       16       17      100
X17     jtl_base_test       17       18      100
X18     jtl_base_test       18       19      100
X19     jtl_base_test       19       20      100
X20     jtl_base_test       20       21      100
.ends
** + -------------------- +

*** top cell: DCHFQ - HFQJTL
Vin1                    1       0       PWL(0ps 0mV   500ps 0mV 501ps 0.517mV 502ps 0.517mV 503ps 0mV  600ps 0mV 601ps 0.517mV 602ps 0.517mV 603ps 0mV)
R1                      1       11      1ohm
X1      jtl_base8       11      12      100        
X2      jtl_base8       12      13      100   
X3      jtl_base8       13      14      100   
X4      jtl_base8       14      15      100 

X35     jtl_base20      15      25      100

X5      jtl_base8       25      26      100        
X6      jtl_base8       26      27      100   
X7      jtl_base8       27      28      100   
X8      jtl_base8       28      76      100   
R72                         76      77 6.592249674902471ohm
L1                      77      0       2pH
Vb1                         100     0                       pwl(0ps 0mV 100ps 0.5mv)

* .tran 0.1ps 1300ps 0ps 0.1ps
.tran 0.1ps 1700ps 0ps 0.1ps

.print phase B1|X1|X1|X35
.print phase B2|X1|X1|X35

.print phase B1|X2|X20|X35
.print phase B2|X2|X20|X35
.print devv  R1

.print phase B1|X1|X2|X2
.print phase B2|X1|X2|X2
.print phase B1|X2|X6|X7
.print phase B2|X2|X6|X7
.print phase B1|X1|X1|X5
.print phase B2|X1|X1|X5
.end